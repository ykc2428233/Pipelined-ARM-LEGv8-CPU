LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SingleCycleCPU_tb IS
END SingleCycleCPU_tb;

ARCHITECTURE tb OF SingleCycleCPU_tb IS
  SIGNAL clk : STD_LOGIC;
  SIGNAL rst : STD_LOGIC;
  SIGNAL DEBUG_PC : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL DEBUG_INSTRUCTION : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL DEBUG_TMP_REGS : STD_LOGIC_VECTOR(64*4 - 1 DOWNTO 0);
  SIGNAL DEBUG_SAVED_REGS : STD_LOGIC_VECTOR(64*4 - 1 DOWNTO 0);
  SIGNAL DEBUG_MEM_CONTENTS : STD_LOGIC_VECTOR(64*4 - 1 DOWNTO 0);
  --SIGNAL TMP_DEBUG : STD_LOGIC_VECTOR(63 DOWNTO 0);
  --SIGNAL TMP_OPcode : STD_LOGIC_VECTOR(3 DOWNTO 0);
  --SIGNAL DEBUG_Reg2Loc : STD_LOGIC;
  --SIGNAL DEBUG_CBranch : STD_LOGIC;
  --SIGNAL DEBUG_MemRead : STD_LOGIC;
  --SIGNAL DEBUG_MemtoReg : STD_LOGIC;
  --SIGNAL DEBUG_MemWrite : STD_LOGIC;
  --SIGNAL DEBUG_ALUSrc : STD_LOGIC;
  --SIGNAL DEBUG_RegWrite : STD_LOGIC;
  --SIGNAL DEBUG_UBranch : STD_LOGIC;
  --SIGNAL DEBUG_ALUOp : STD_LOGIC_VECTOR(1 DOWNTO 0);
  --SIGNAL DEBUG_ZERO : STD_LOGIC;

BEGIN
  UUT_CPU : ENTITY work.SingleCycleCPU	
    PORT MAP(
	clk => clk,
	rst => rst,
	DEBUG_PC => DEBUG_PC,
	DEBUG_TMP_REGS => DEBUG_TMP_REGS,
	DEBUG_SAVED_REGS => DEBUG_SAVED_REGS,
	DEBUG_MEM_CONTENTS => DEBUG_MEM_CONTENTS,
        DEBUG_INSTRUCTION => DEBUG_INSTRUCTION
        --TMP_DEBUG => TMP_DEBUG,
	--TMP_OPcode => TMP_OPcode,
	--DEBUG_Reg2Loc => DEBUG_Reg2Loc,
  	--DEBUG_CBranch => DEBUG_CBranch,
  	--DEBUG_MemRead => DEBUG_MemRead,
  	--DEBUG_MemtoReg => DEBUG_MemtoReg,
 	--DEBUG_MemWrite => DEBUG_MemWrite,
 	--DEBUG_ALUSrc => DEBUG_ALUSrc,
  	--DEBUG_RegWrite => DEBUG_RegWrite,
 	--DEBUG_UBranch => DEBUG_UBranch,
 	--DEBUG_ALUOp => DEBUG_ALUOp,
	--DEBUG_ZERO => DEBUG_ZERO
    );
  
  clock : PROCESS
    CONSTANT clk_period : TIME := 50 ns;
    BEGIN
      clk <= '1';
      WAIT FOR clk_period;
      clk <= '0';
      WAIT FOR clk_period;
    END PROCESS;

  reset : PROCESS
    BEGIN
      rst <= '1';
      WAIT FOR 10 ns;
      rst <= '0';
      WAIT FOR 100 ms;
    END PROCESS;

END tb;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
 
ENTITY EQUAL0 IS
PORT(
	datavalue : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
	eq0 : OUT STD_LOGIC
    );
END EQUAL0;

ARCHITECTURE behavioral of EQUAL0 IS
CONSTANT ZR : STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS => '0');
BEGIN
  PROCESS(datavalue)
  BEGIN
  IF (datavalue(63 DOWNTO 0) = x"0000000000000000") THEN
    eq0 <= '1';
  ELSE
    eq0 <= '0';
  END IF;
  END PROCESS;

END behavioral;
